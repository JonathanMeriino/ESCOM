Cypress C22V10 Jedec Fuse File: led.jed

This file was created on 03/28/2021 at 20:18:55 
by PLA2JED.EXE    31/03/2000  [v4.02 ] 6.3 IR 35

C22V10*
QP24*                Number of Pins*
QF5828*              Number of Fuses*
F0*                  Note: Default fuse setting 0*
G0*                  Note: Security bit Unprogrammed*
NOTE DEVICE C22V10*
NOTE PACKAGE palce22v10-25pc/pi*
NOTE PROPERTY BUS_HOLD ENABLE*
NOTE PINS  a(4):1 a(3):2 a(2):3 a(1):4 a(0):5 sal(4):14 sal(2):15 sal(0):16 *
NOTE PINS  sal(1):22 sal(3):23 *
NOTE PINS *
NOTE NODES *
L00000
00000000000000000000000000000000000000000000
* Node a(4)[1] => BANK : 1 *

L00044
11111111111111111111111111111111111111111111
11110111111111111111111111111111111111111111
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
* Node sal(3)[23] => OE : 1 ,LOGIC : 8 *

L00440
11111111111111111111111111111111111111111111
11111111111101111111111111111111111111111111
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
* Node sal(1)[22] => OE : 1 ,LOGIC : 10 *

L00924
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
* Not Used #[21] => OE : 1 ,LOGIC : 12 *

L01496
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
* Not Used #[20] => OE : 1 ,LOGIC : 14 *

L02156
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
* Not Used #[19] => OE : 1 ,LOGIC : 16 *

L02904
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
* Not Used #[18] => OE : 1 ,LOGIC : 16 *

L03652
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
* Not Used #[17] => OE : 1 ,LOGIC : 14 *

L04312
11111111111111111111111111111111111111111111
11111111111111110111111111111111111111111111
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
* Node sal(0)[16] => OE : 1 ,LOGIC : 12 *

L04884
11111111111111111111111111111111111111111111
11111111011111111111111111111111111111111111
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
* Node sal(2)[15] => OE : 1 ,LOGIC : 10 *

L05368
11111111111111111111111111111111111111111111
01111111111111111111111111111111111111111111
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000
* Node sal(4)[14] => OE : 1 ,LOGIC : 8 *

L05764
00000000000000000000000000000000000000000000
* Node a(3)[2] => BANK : 1 *

L05808
11* Note: 23 *

L05810
11* Note: 22 *

L05812
00* Note: 21 *

L05814
00* Note: 20 *

L05816
00* Note: 19 *

L05818
00* Note: 18 *

L05820
00* Note: 17 *

L05822
11* Note: 16 *

L05824
11* Note: 15 *

L05826
11* Note: 14 *

C3775*               Note: Fuse Checksum*
6E26
